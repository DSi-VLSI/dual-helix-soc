module dummy_rtl;

  initial begin
    $display("This is a dummy RTL module.");
  end

endmodule
