package soc_ctrl_pkg;

  parameter int REF_DIV_BW = 4;
  parameter int FB_DIV_BW = 12;

endpackage
